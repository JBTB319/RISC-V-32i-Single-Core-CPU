hdl/components/alu.sv
hdl/components/data_memory.sv
hdl/components/instruction_memory.sv
hdl/components/program_counter.sv
hdl/components/register_file.sv
hdl/components/sign_extender.sv

