module tb_instruction_memory;

endmodule