module alu (
   input logic [31:0] srcA,
   input logic [31:0] srcB,
   input logic [2:0] aluSel,
   output logic [31:0] aluResult
);

endmodule